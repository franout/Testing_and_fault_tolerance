LIBRARY ieee;
USE ieee.std_logic_1164.ALL;


ENTITY  circ4 IS
PORT ( clk, reset, cnt: IN std_logic;
		y: OUT std_logic);
END ENTITY circ4;

ARCHITECTURE struc OF circ4 IS


BEGIN






regs:PROCESS()
BEGIN 

END PROCESS regs;



logic:PROCESS()
BEGIN


END PROCESS logic;

END struc;
